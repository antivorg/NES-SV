/*
*
* ALU
*
*/

module ALU (
    input logic [7:0] A, B,
    input logic statusReg[7:0],
    input logic decEnable, carrIn,
    output logic [7:0] resultReg,
    output logic overFlow, carrOut, halfCarry, 
);

    

endmodule