/*
*   Data Bus
*/

interface dataBus;
    wire A[15:0];
    wire D[7:0];
    logic write;
endinterface